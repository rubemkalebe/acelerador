library ieee;
use ieee.std_logic_1164.all;

entity basic_unit is
  generic (
    n : natural := 32
  );
end basic_unit;

architecture basic_unit of basic_unit is

  signal

begin

end basic_unit;
