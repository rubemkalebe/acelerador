-- Short description...
-- Version: 03.08.2016.

library ieee;
use ieee.std_logic_1164.all;

entity load_store is
end load_store;

architecture load_store of load_store is

begin
  
end load_store;
