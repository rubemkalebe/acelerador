library ieee;
use ieee.std_logic_1164.all;

entity accelerator is
  generic (
    n : natural := 32
  );
end accelerator;

architecture accelerator of accelerator is

  signal

begin

end accelerator;
