library ieee;
use ieee.std_logic_1164.all;

entity cluster is
  generic (
    n : natural := 32
  );
end cluster;

architecture cluster of cluster is

  signal

begin

end cluster;
