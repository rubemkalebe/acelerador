library ieee;
use ieee.std_logic_1164.all;

entity register_file is
  generic (
    n : natural := 32
  );
end register_file;

architecture register_file of register_file is

  signal

begin

end register_file;
