library ieee;
use ieee.std_logic_1164.all;

entity global_register_file is
  generic (
    n : natural := 32
  );
end global_register_file;

architecture global_register_file of global_register_file is

  signal

begin

end global_register_file;
